`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// 基本完成 
// 
//////////////////////////////////////////////////////////////////////////////////
module ID(clk,Instruction_id, PC_id, RegWrite_wb, rdAddr_wb, RegWriteData_wb, MemRead_ex, 
          rdAddr_ex, MemtoReg_id, RegWrite_id, MemWrite_id, MemRead_id, ALUCode_id, 
			 ALUSrcA_id, ALUSrcB_id,  Stall, Branch, Jump, IFWrite,  JumpAddr, Imm_id,
			 rs1Data_id, rs2Data_id,rs1Addr_id,rs2Addr_id,rdAddr_id);
    input clk;
    input [31:0] Instruction_id;
    input [31:0] PC_id;
    input RegWrite_wb;
    input [4:0] rdAddr_wb;
    input [31:0] RegWriteData_wb;
    input MemRead_ex;
    input [4:0] rdAddr_ex;
    output MemtoReg_id;
    output RegWrite_id;
    output MemWrite_id;
    output MemRead_id;
    output [3:0] ALUCode_id;
    output ALUSrcA_id;
    output [1:0]ALUSrcB_id;
    output Stall;
    output Branch;
    output Jump;
    output IFWrite;
    output [31:0] JumpAddr;
    output [31:0] Imm_id;
    output [31:0] rs1Data_id;
    output [31:0] rs2Data_id;
	output[4:0] rs1Addr_id,rs2Addr_id,rdAddr_id;

    wire [31:0] offset;
    wire JALR;
    wire [31:0] JALR_Addr;
 
    // Decode
    Decode Decode1(
        .Instruction(Instruction_id),	// current instruction
        .MemtoReg(MemtoReg_id),		// use memory output as into register
        .RegWrite(RegWrite_id),		// enable writing back to 
        .MemWrite(MemWrite_id),		// write to memory
        .MemRead(MemRead_id),
        .ALUCode(ALUCode_id),         // ALU operation select
        .ALUSrcA(ALUSrcA_id),
        .ALUSrcB(ALUSrcB_id),
        .Jump(JUMP),
        .JALR(JALR),
        .Imm(Imm_id),
        .offset(offset)
    );


    // Registers 
    Registers Registers1(
        .clk(clk), 
        .rs1Addr(rs1Addr_id), 
        .rs2Addr(rs2Addr_id), 
        .WriteAddr(rdAddr_wb), 
        .RegWrite(RegWrite_wb), 
        .WriteData(RegWriteData_wb), 
        .rs1Data(rs1Data_id), 
        .rs2Data(rs2Data_id)
    ); 

    // Hazard Detector
    assign Stall = ((rdAddr_ex == rs1Addr_id)||(rdAddr_ex == rs2Addr_id))&&MemRead_ex;
    assign IFWrite = ~Stall;

    // BranchTest 
    BranchTest BranchTest1(
        .Instruction(Instruction_id), 
        .rs1Data(rs1Data_id), 
        .rs2Data(rs2Data_id), 
        .Branch(Branch)
    );


    // 二路选择器
    mux_2to1 mux1(
        .addr(JALR),
        .in0(PC_id),
        .in1(rs1Data_id),
        .out(JALR_Addr)
    );
    adder_32bits addr32(
        .a(JALR_Addr),
        .b(offset),
        .ci(0),
        .s(JumpAddr),
        .co()
    );
    
endmodule

module BranchTest (
    ports
);
    
endmodule